    Mac OS X            	   2        2                                      ATTR      2   �   v                  �   #  com.apple.quarantine    �   S  com.dropbox.attributes   q/0002;554e1bda;The\x20Unarchiver; x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK���lK}�J� ��"����|_S�t[[���Z ���