-- ====================================================================
--
--	File Name:		Test_Counter.vhd
--	Description:	Test bench for counter 
--					
--
--	Date:			15/03/2013
--	Designer:		Amiram Lifshitz & Amit Biran
--		
-- ====================================================================
-- MIPS PIPELINE Stage I - Instruction Fetch.			

LIBRARY IEEE; 			
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;